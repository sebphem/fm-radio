module demodulate #(
    parameter DATA_WIDTH=32
) (
    input logic [(DATA_WIDTH-1):0] real;
    input logic [(DATA_WIDTH1):0] imag;
    input logic [(DATA_WIDTH1):0] real_prev;
    input logic [(DATA_WIDTH-1):0] real;
);
    
endmodule