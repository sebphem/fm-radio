package synth_global


    localparam BITS = 10
    localparam QUANT_VAL = (1 << BITS);

    function int QUANTIZE_I(int i);
        return i * QUANT_VAL;
    endfunction


    function int DEQUANTIZE_I(int i);
        return i / QUANT_VAL;
    endfunction
    localparam AUDIO_DECIM = 8;
    localparam SAMPLES = 65536*4;
    localparam AUDIO_SAMPLES = SAMPLES/AUDIO_DECIM;
    localparam MAX_TAPS = 32;

    logic [31:0] channel_coeffs_real [19:0] = '{
        32'h00000001, 32'h00000008, 32'hfffffff3, 32'h00000009, 
        32'h0000000b, 32'hffffffd3, 32'h00000045, 32'hffffffd3, 
        32'hffffffb1, 32'h00000257, 32'h00000257, 32'hffffffb1, 
        32'hffffffd3, 32'h00000045, 32'hffffffd3, 32'h0000000b, 
        32'h00000009, 32'hfffffff3, 32'h00000008, 32'h00000001
    };

    logic [31:0] channel_coeffs_imag [19:0] = '{
        32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
        32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
        32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
        32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
        32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
    };

    localparam int AUDIO_LPR_COEFF_TAPS = 32;
    logic [31:0] audio_lpr_coeffs [31:0] = '{
        32'hfffffffd, 32'hfffffffa, 32'hfffffff4, 32'hffffffed, 
        32'hffffffe5, 32'hffffffdf, 32'hffffffe2, 32'hfffffff3, 
        32'h00000015, 32'h0000004e, 32'h0000009b, 32'h000000f9, 
        32'h0000015d, 32'h000001be, 32'h0000020e, 32'h00000243, 
        32'h00000243, 32'h0000020e, 32'h000001be, 32'h0000015d, 
        32'h000000f9, 32'h0000009b, 32'h0000004e, 32'h00000015, 
        32'hfffffff3, 32'hffffffe2, 32'hffffffdf, 32'hffffffe5, 
        32'hffffffed, 32'hfffffff4, 32'hfffffffa, 32'hfffffffd
    };

    localparam int AUDIO_LMR_COEFF_TAPS = 32;
    logic [31:0] audio_lmr_coeffs [31:0] = '{
        32'hfffffffd, 32'hfffffffa, 32'hfffffff4, 32'hffffffed, 
        32'hffffffe5, 32'hffffffdf, 32'hffffffe2, 32'hfffffff3, 
        32'h00000015, 32'h0000004e, 32'h0000009b, 32'h000000f9, 
        32'h0000015d, 32'h000001be, 32'h0000020e, 32'h00000243, 
        32'h00000243, 32'h0000020e, 32'h000001be, 32'h0000015d, 
        32'h000000f9, 32'h0000009b, 32'h0000004e, 32'h00000015, 
        32'hfffffff3, 32'hffffffe2, 32'hffffffdf, 32'hffffffe5, 
        32'hffffffed, 32'hfffffff4, 32'hfffffffa, 32'hfffffffd
    };

    localparam int BP_PILOT_COEFF_TAPS = 32;
    logic [31:0] bp_pilot_coeffs [31:0] = '{
        32'h0000000e, 32'h0000001f, 32'h00000034, 32'h00000048, 
        32'h0000004e, 32'h00000036, 32'hfffffff8, 32'hffffff98, 
        32'hffffff2d, 32'hfffffeda, 32'hfffffec3, 32'hfffffefe, 
        32'hffffff8a, 32'h0000004a, 32'h0000010f, 32'h000001a1, 
        32'h000001a1, 32'h0000010f, 32'h0000004a, 32'hffffff8a, 
        32'hfffffefe, 32'hfffffec3, 32'hfffffeda, 32'hffffff2d, 
        32'hffffff98, 32'hfffffff8, 32'h00000036, 32'h0000004e, 
        32'h00000048, 32'h00000034, 32'h0000001f, 32'h0000000e
    };

    localparam int BP_LMR_COEFF_TAPS = 32;
    logic [31:0] bp_lmr_coeffs [31:0] = '{
        32'h00000000, 32'h00000000, 32'hfffffffc, 32'hfffffff9, 
        32'hfffffffe, 32'h00000008, 32'h0000000c, 32'h00000002, 
        32'h00000003, 32'h0000001e, 32'h00000030, 32'hfffffffc, 
        32'hffffff8c, 32'hffffff58, 32'hffffffc3, 32'h0000008a, 
        32'h0000008a, 32'hffffffc3, 32'hffffff58, 32'hffffff8c, 
        32'hfffffffc, 32'h00000030, 32'h0000001e, 32'h00000003, 
        32'h00000002, 32'h0000000c, 32'h00000008, 32'hfffffffe, 
        32'hfffffff9, 32'hfffffffc, 32'h00000000, 32'h00000000
    };

    localparam int HP_COEFF_TAPS = 32;
    logic [31:0] hp_coeffs [31:0] = '{
        32'hffffffff, 32'h00000000, 32'h00000000, 32'h00000002, 
        32'h00000004, 32'h00000008, 32'h0000000b, 32'h0000000c, 
        32'h00000008, 32'hffffffff, 32'hffffffee, 32'hffffffd7, 
        32'hffffffbb, 32'hffffff9f, 32'hffffff87, 32'hffffff76, 
        32'hffffff76, 32'hffffff87, 32'hffffff9f, 32'hffffffbb, 
        32'hffffffd7, 32'hffffffee, 32'hffffffff, 32'h00000008, 
        32'h0000000c, 32'h0000000b, 32'h00000008, 32'h00000004, 
        32'h00000002, 32'h00000000, 32'h00000000, 32'hffffffff
    };

    logic [31:0] sin_lut [1023:0] = '{
        32'h00000000, 32'h00000006, 32'h0000000C, 32'h00000012, 32'h00000019, 32'h0000001F, 32'h00000025, 32'h0000002B, 
        32'h00000032, 32'h00000038, 32'h0000003E, 32'h00000045, 32'h0000004B, 32'h00000051, 32'h00000057, 32'h0000005E, 
        32'h00000064, 32'h0000006A, 32'h00000070, 32'h00000077, 32'h0000007D, 32'h00000083, 32'h00000089, 32'h00000090, 
        32'h00000096, 32'h0000009C, 32'h000000A2, 32'h000000A8, 32'h000000AF, 32'h000000B5, 32'h000000BB, 32'h000000C1, 
        32'h000000C7, 32'h000000CD, 32'h000000D4, 32'h000000DA, 32'h000000E0, 32'h000000E6, 32'h000000EC, 32'h000000F2, 
        32'h000000F8, 32'h000000FE, 32'h00000104, 32'h0000010B, 32'h00000111, 32'h00000117, 32'h0000011D, 32'h00000123, 
        32'h00000129, 32'h0000012F, 32'h00000135, 32'h0000013B, 32'h00000141, 32'h00000147, 32'h0000014D, 32'h00000153, 
        32'h00000158, 32'h0000015E, 32'h00000164, 32'h0000016A, 32'h00000170, 32'h00000176, 32'h0000017C, 32'h00000182, 
        32'h00000187, 32'h0000018D, 32'h00000193, 32'h00000199, 32'h0000019E, 32'h000001A4, 32'h000001AA, 32'h000001B0, 
        32'h000001B5, 32'h000001BB, 32'h000001C1, 32'h000001C6, 32'h000001CC, 32'h000001D2, 32'h000001D7, 32'h000001DD, 
        32'h000001E2, 32'h000001E8, 32'h000001ED, 32'h000001F3, 32'h000001F8, 32'h000001FE, 32'h00000203, 32'h00000209, 
        32'h0000020E, 32'h00000213, 32'h00000219, 32'h0000021E, 32'h00000223, 32'h00000229, 32'h0000022E, 32'h00000233, 
        32'h00000238, 32'h0000023E, 32'h00000243, 32'h00000248, 32'h0000024D, 32'h00000252, 32'h00000257, 32'h0000025C, 
        32'h00000261, 32'h00000267, 32'h0000026C, 32'h00000271, 32'h00000275, 32'h0000027A, 32'h0000027F, 32'h00000284, 
        32'h00000289, 32'h0000028E, 32'h00000293, 32'h00000298, 32'h0000029C, 32'h000002A1, 32'h000002A6, 32'h000002AB, 
        32'h000002AF, 32'h000002B4, 32'h000002B8, 32'h000002BD, 32'h000002C2, 32'h000002C6, 32'h000002CB, 32'h000002CF, 
        32'h000002D4, 32'h000002D8, 32'h000002DC, 32'h000002E1, 32'h000002E5, 32'h000002E9, 32'h000002EE, 32'h000002F2, 
        32'h000002F6, 32'h000002FA, 32'h000002FF, 32'h00000303, 32'h00000307, 32'h0000030B, 32'h0000030F, 32'h00000313, 
        32'h00000317, 32'h0000031B, 32'h0000031F, 32'h00000323, 32'h00000327, 32'h0000032B, 32'h0000032E, 32'h00000332, 
        32'h00000336, 32'h0000033A, 32'h0000033D, 32'h00000341, 32'h00000345, 32'h00000348, 32'h0000034C, 32'h0000034F, 
        32'h00000353, 32'h00000356, 32'h0000035A, 32'h0000035D, 32'h00000361, 32'h00000364, 32'h00000367, 32'h0000036B, 
        32'h0000036E, 32'h00000371, 32'h00000374, 32'h00000377, 32'h0000037A, 32'h0000037E, 32'h00000381, 32'h00000384, 
        32'h00000387, 32'h0000038A, 32'h0000038C, 32'h0000038F, 32'h00000392, 32'h00000395, 32'h00000398, 32'h0000039A, 
        32'h0000039D, 32'h000003A0, 32'h000003A2, 32'h000003A5, 32'h000003A8, 32'h000003AA, 32'h000003AD, 32'h000003AF, 
        32'h000003B2, 32'h000003B4, 32'h000003B6, 32'h000003B9, 32'h000003BB, 32'h000003BD, 32'h000003BF, 32'h000003C2, 
        32'h000003C4, 32'h000003C6, 32'h000003C8, 32'h000003CA, 32'h000003CC, 32'h000003CE, 32'h000003D0, 32'h000003D2, 
        32'h000003D3, 32'h000003D5, 32'h000003D7, 32'h000003D9, 32'h000003DA, 32'h000003DC, 32'h000003DE, 32'h000003DF, 
        32'h000003E1, 32'h000003E2, 32'h000003E4, 32'h000003E5, 32'h000003E7, 32'h000003E8, 32'h000003E9, 32'h000003EB, 
        32'h000003EC, 32'h000003ED, 32'h000003EE, 32'h000003EF, 32'h000003F0, 32'h000003F1, 32'h000003F2, 32'h000003F3, 
        32'h000003F4, 32'h000003F5, 32'h000003F6, 32'h000003F7, 32'h000003F8, 32'h000003F9, 32'h000003F9, 32'h000003FA, 
        32'h000003FB, 32'h000003FB, 32'h000003FC, 32'h000003FC, 32'h000003FD, 32'h000003FD, 32'h000003FE, 32'h000003FE, 
        32'h000003FE, 32'h000003FF, 32'h000003FF, 32'h000003FF
    };


endpackage