package synth_func
    
    function int QUANTIZE_I(int i);
        return i * QUANT_VAL;
    endfunction
 
endpackage