module iir #(
    parameter DATA_WIDTH = 32;
    
) (
    ports
);
    
endmodule